package pkg_verification
  `include "cls_dump_ctrl_f.sv"
  `include "cls_dump_ctrl_l.sv"
  `include "cls_dump_ppm.sv"
endpackage

