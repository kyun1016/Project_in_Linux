// 
`define DIR_TB_TOP u_tb_top
`define DIR_TX_TOP `DIR_TB_TOP.u_tx_top

