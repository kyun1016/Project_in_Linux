package pkg_tx_data;
  `include "cls_clock_train_pattern.sv"
  `include "cls_ctrl_f.sv"
  `include "cls_ctrl_l.sv"
//   `include "cls_image.sv"
  `include "cls_k_symbol.sv"
  `include "cls_link_stable_pattern.sv"
endpackage

