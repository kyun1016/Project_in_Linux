// ../../list_tx_model.f

package pkg_tx_sequencer;
  `include "cls_sequencer.sv"
endpackage

